module EXP_GATE_2(input A,input B,input C,output X); // This is IC 7462
assign X = A & B & C;
endmodule
